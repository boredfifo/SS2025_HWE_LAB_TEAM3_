ENTITY ALU_DECODER IS
PORT(F0, F1: IN BIT;
	F_00, F_01, F_10, F_11: OUT BIT);
END ALU_DECODER;

ARCHITECTURE behavioural of ALU_DECODER IS
SIGNAL F0_NOT, F1_NOT: BIT;

BEGIN

F0_NOT<= NOT F0;
F1_NOT<= NOT F1;

F_00<=	F0_NOT AND F1_NOT;
F_01<=	F0_NOT AND F1;
F_10<=	F0 AND F1_NOT;
F_11<=	F0 and F1;

END behavioural;
